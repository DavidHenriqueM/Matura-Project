`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.06.2023 12:22:38
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// state maschine that interprets commands

module top(
    input sys_clk,
    input sw_0, // reset
    input RsRx,
    output RsTx
    );

    
    wire         mem_readWrite;
    wire [31:0]  mem_dataIn;
    wire         mem_enable;
    wire [14:0]   mem_address;
    wire [31:0] mem_dataOut;

    //registers and wires for memory arbitrator

    reg memJudge_enable = 1;
    wire Judge_mem_enable1;
    wire Judge_mem_enable2;
    wire Judge_mem_readWrite1;
    wire Judge_mem_readWrite2; 
    wire [14:0] Judge_Address1;
    wire [14:0] Judge_Address2;
    wire [31:0] Judge_data1;
    wire [31:0] Judge_data2;
    wire [31:0] Judge_DataOut1;
    wire [31:0] Judge_DataOut2;
    wire Judge_done1;
    wire Judge_done2;

    wire        exec_done;
    wire [31:0] exec_data;
    wire        exec_sample;

    TopUART TopUART(
       .clk             (sys_clk),
       .rst             (sw_0),
       .serial_in       (RsRx),
       .arbitratorDone  (Judge_done1),
       .dataOutOfMemory (Judge_DataOut1), 
       .serial_out      (RsTx),
       .out_readWrite   (Judge_mem_readWrite1),
       .dataIntoMemory  (Judge_data1),
       .memoryEnable    (Judge_mem_enable1),
       .memoryAddress   (Judge_Address1)
    );


    memoryArbitration memJudge(
        .clock         (sys_clk),
        .reset         (sw_0),
        .moduleEnable  (memJudge_enable),
        .memoryEnable1 (Judge_mem_enable1),
        .memoryEnable2 (Judge_mem_enable2),
        .readWrite1    (Judge_mem_readWrite1),
        .readWrite2    (Judge_mem_readWrite2),
        .Address1      (Judge_Address1),
        .Address2      (Judge_Address2),
        .Data1         (Judge_data1),
        .Data2         (Judge_data2),
        .DataOut1      (Judge_DataOut1),
        .DataOut2      (Judge_DataOut2),
        .done1         (Judge_done1),
        .done2         (Judge_done2)
        );

    ringBuffer ringBuffer(
        .clk               (sys_clk),
        .rst               (sw_0),
        .mem_DataOut       (Judge_DataOut2),
        .mem_done          (Judge_done2),
        .exec_done         (exec_done),
        .mem_enable        (Judge_mem_enable2),
        .mem_readWrite     (Judge_mem_readWrite2),
        .mem_address       (Judge_Address2),
        .mem_DataWrite     (Judge_data2),
        .dataToInterpreter (exec_data),
        .exec_sample       (exec_sample)
        );

endmodule