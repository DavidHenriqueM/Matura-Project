`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/13/2023 09:01:27 AM
// Design Name: 
// Module Name: seq_to_matrix
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module seq_to_matrix(
    input clock,
    input reset,
    input [31:0]data_In,
    input sizeX,
    input sizeY,
    output reg [31:0] out_Matrix [0:31][0:31],
    output reg done
    );





endmodule
